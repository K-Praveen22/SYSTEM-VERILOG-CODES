// Code your design here
module add(input [3:0]a,
           input [3:0]b,
           output [5:0]c );
  assign c =a+b;
endmodule
    
